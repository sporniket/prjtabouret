module top(i2, i3, m1);

input i2;
input i3;
output m1;

assign m1 = i2 & i3;
endmodule
